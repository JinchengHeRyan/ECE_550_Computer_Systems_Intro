module add_circuit(result, data_A, data_B);
  output [31:0] result;
  input [31:0] data_A;
  input [31:0] data_B;


endmodule
